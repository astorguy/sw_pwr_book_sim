** Sheet_1 **
VEASYEDA EASYEDA GND 1
RUPPER DIV OUT 10K
RLOWER VEE DIV 10K
E1 Q1_BASE VEE VEE DIV 10K
Q1 OUT Q1_BASE IN 2N2222

.tran 1m 3.1415
.inc standard.bjt

** Sheet_1 **
VEASYEDA EASYEDA GND 1
R1 IN OUT1 140
R2 IN OUT2 132
.TRAN 1M 3.1415

** Sheet_1 **
VEASYEDA EASYEDA GND 1
R1 IN MID 1K
C1 COM MID 0.1U
R2 MID OUT 100
.tran 1m 3.1415

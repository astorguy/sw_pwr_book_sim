.title KiCad schematic
E2 base vee ref div 10k
Q1 in base out 2N2222   
RLOWER1 div vee 100
RUPPER1 out div 50
.end

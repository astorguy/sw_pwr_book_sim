** Sheet_1 **
VEASYEDA EASYEDA GND 1
R1 IN OUT1 140
R2 IN OUT2 132
.tran 1m 3.1415

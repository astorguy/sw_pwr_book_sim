* title line

rlower1 div com 10k
e1 beta com vref div 100
rupper1 out div 10k
e2 g com beta com 10
x2 in gain gain k=0.05
rsol1 sum out 1
x3 gain g sum sum k1=1 k2=1 a=1
rf rc beta 100
cf rc div 100n
iload out 0 ac 1

vcom com 0 dc 0
vref vref 0 dc 2.5

vin in 0 dc 15

.subckt gain in out k=1
e1 out 0 in 0 {k}
.ends gain

.subckt sum in1 in2 out k1=1 k2=1 a=1
b1 out 0 v = {a * ((v(in1) * k1) + (v(in2) * k2))}
.ends sum

.control
* timestamp: tue apr  2 22:38:22 2024
set wr_singlescale  $ makes one x-axis for wrdata
set wr_vecnames     $ puts names at top of columns
ac dec 100 10m 100k
wrdata /workspaces/sw_pwr_book_sim/circuits/sec_1_04_04_lin_reg/sim_results/ac1.txt 20*log10(mag(out))
quit
.endc
.end